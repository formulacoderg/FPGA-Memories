module tb_rtl_crack();

// Your testbench goes here.

endmodule: tb_rtl_crack
