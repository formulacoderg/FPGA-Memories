module tb_rtl_task4();

// Your testbench goes here.

endmodule: tb_rtl_task4
